-- jtag_uart.vhd

-- Generated using ACDS version 20.1 720


package jtag_uart1 is
component jtag_uart is
	port (
		avalon_jtag_slave_chipselect  : in  std_logic                     := '0';             -- avalon_jtag_slave.chipselect
		avalon_jtag_slave_address     : in  std_logic                     := '0';             --                  .address
		avalon_jtag_slave_read_n      : in  std_logic                     := '0';             --                  .read_n
		avalon_jtag_slave_readdata    : out std_logic_vector(31 downto 0);                    --                  .readdata
		avalon_jtag_slave_write_n     : in  std_logic                     := '0';             --                  .write_n
		avalon_jtag_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		avalon_jtag_slave_waitrequest : out std_logic;                                        --                  .waitrequest
		clk_1_clk                     : in  std_logic                     := '0';             --             clk_1.clk
		irq_irq                       : out std_logic;                                        --               irq.irq
		reset_1_reset_n               : in  std_logic                     := '0'              --           reset_1.reset_n
	);
end component jtag_uart;
end package jtag_uart1;

--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.numeric_std.all;

entity jtag_uart is
	port (
		avalon_jtag_slave_chipselect  : in  std_logic                     := '0';             -- avalon_jtag_slave.chipselect
		avalon_jtag_slave_address     : in  std_logic                     := '0';             --                  .address
		avalon_jtag_slave_read_n      : in  std_logic                     := '0';             --                  .read_n
		avalon_jtag_slave_readdata    : out std_logic_vector(31 downto 0);                    --                  .readdata
		avalon_jtag_slave_write_n     : in  std_logic                     := '0';             --                  .write_n
		avalon_jtag_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		avalon_jtag_slave_waitrequest : out std_logic;                                        --                  .waitrequest
		clk_1_clk                     : in  std_logic                     := '0';             --             clk_1.clk
		irq_irq                       : out std_logic;                                        --               irq.irq
		reset_1_reset_n               : in  std_logic                     := '0'              --           reset_1.reset_n
	);
end entity jtag_uart;

architecture rtl of jtag_uart is
	component jtag_uart_ju is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component jtag_uart_ju;

begin

	ju : component jtag_uart_ju
		port map (
			clk            => clk_1_clk,                     --               clk.clk
			rst_n          => reset_1_reset_n,               --             reset.reset_n
			av_chipselect  => avalon_jtag_slave_chipselect,  -- avalon_jtag_slave.chipselect
			av_address     => avalon_jtag_slave_address,     --                  .address
			av_read_n      => avalon_jtag_slave_read_n,      --                  .read_n
			av_readdata    => avalon_jtag_slave_readdata,    --                  .readdata
			av_write_n     => avalon_jtag_slave_write_n,     --                  .write_n
			av_writedata   => avalon_jtag_slave_writedata,   --                  .writedata
			av_waitrequest => avalon_jtag_slave_waitrequest, --                  .waitrequest
			av_irq         => irq_irq                        --               irq.irq
		);

end architecture rtl; -- of jtag_uart
